LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;
USE work.aux_package.all;
------------------------------------------------------------------
entity segment is
	generic ( n : positive := 8 ); 
	port(num1 : in std_logic_vector(3 downto 0);
		 num2: in std_logic_vector(3 downto 0);
		 out_h1 : out std_logic_vector(6 downto 0);
		 out_h2 : out std_logic_vector(6 downto 0));
end segment;
------------------------------------------------------------------
architecture arc_sys of segment is	
SIGNAL NUM_e1 : integer ;
SIGNAL NUM_e2 : integer ;
begin
    
	with num1 select
		out_h1<=(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'0',6=>'1') when "0000",
				(0=>'1',1=>'0',2=>'0',3=>'1',4=>'1',5=>'1',6=>'1') when "0001",
				(0=>'0',1=>'0',2=>'1',3=>'0',4=>'0',5=>'1',6=>'0') when "0010",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'1',5=>'1',6=>'0') when "0011",
				(0=>'1',1=>'0',2=>'0',3=>'1',4=>'1',5=>'0',6=>'0') when "0100",
				(0=>'0',1=>'1',2=>'0',3=>'0',4=>'1',5=>'0',6=>'0') when "0101",
				(0=>'0',1=>'1',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "0110",
				(0=>'0',1=>'0',2=>'0',3=>'1',4=>'1',5=>'1',6=>'1') when "0111",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "1000",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'1',5=>'0',6=>'0') when "1001",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'1',6=>'0') when "1010",
				(0=>'1',1=>'1',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "1011",
				(0=>'0',1=>'1',2=>'1',3=>'0',4=>'0',5=>'0',6=>'1') when "1100",
				(0=>'1',1=>'0',2=>'0',3=>'0',4=>'0',5=>'1',6=>'0') when "1101",
				(0=>'0',1=>'1',2=>'1',3=>'0',4=>'0',5=>'0',6=>'0') when "1110",
				(0=>'0',1=>'1',2=>'1',3=>'1',4=>'0',5=>'0',6=>'0') when "1111",
				(0=>'1',1=>'1',2=>'1',3=>'1',4=>'1',5=>'1',6=>'1') when others;


	with num2 select
		out_h2<=(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'0',6=>'1') when "0000",
				(0=>'1',1=>'0',2=>'0',3=>'1',4=>'1',5=>'1',6=>'1') when "0001",
				(0=>'0',1=>'0',2=>'1',3=>'0',4=>'0',5=>'1',6=>'0') when "0010",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'1',5=>'1',6=>'0') when "0011",
				(0=>'1',1=>'0',2=>'0',3=>'1',4=>'1',5=>'0',6=>'0') when "0100",
				(0=>'0',1=>'1',2=>'0',3=>'0',4=>'1',5=>'0',6=>'0') when "0101",
				(0=>'0',1=>'1',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "0110",
				(0=>'0',1=>'0',2=>'0',3=>'1',4=>'1',5=>'1',6=>'1') when "0111",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "1000",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'1',5=>'0',6=>'0') when "1001",
				(0=>'0',1=>'0',2=>'0',3=>'0',4=>'0',5=>'1',6=>'0') when "1010",
				(0=>'1',1=>'1',2=>'0',3=>'0',4=>'0',5=>'0',6=>'0') when "1011",
				(0=>'0',1=>'1',2=>'1',3=>'0',4=>'0',5=>'0',6=>'1') when "1100",
				(0=>'1',1=>'0',2=>'0',3=>'0',4=>'0',5=>'1',6=>'0') when "1101",
				(0=>'0',1=>'1',2=>'1',3=>'0',4=>'0',5=>'0',6=>'0') when "1110",
				(0=>'0',1=>'1',2=>'1',3=>'1',4=>'0',5=>'0',6=>'0') when "1111",
				(0=>'1',1=>'1',2=>'1',3=>'1',4=>'1',5=>'1',6=>'1') when others;

end arc_sys;







